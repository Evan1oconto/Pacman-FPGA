library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity ghost_sprite is
  port(
		clk: in std_logic;
		addr : in std_logic_vector(7 downto 0);
		data : out std_logic
  );
end ghost_sprite;



architecture synth of ghost_sprite is
begin
	process(clk) is begin
		if rising_edge(clk) then
			case addr is
			when "00000000" => data <= '0';
			when "00000001" => data <= '0';
			when "00000010" => data <= '0';
			when "00000011" => data <= '0';
			when "00000100" => data <= '0';
			when "00000101" => data <= '0';
			when "00000110" => data <= '0';
			when "00000111" => data <= '0';
			when "00001000" => data <= '0';
			when "00001001" => data <= '0';
			when "00001010" => data <= '0';
			when "00001011" => data <= '0';
			when "00001100" => data <= '0';
			when "00001101" => data <= '0';
			when "00001110" => data <= '0';
			when "00001111" => data <= '0';
			when "00010000" => data <= '0';
			when "00010001" => data <= '0';
			when "00010010" => data <= '0';
			when "00010011" => data <= '0';
			when "00010100" => data <= '0';
			when "00010101" => data <= '0';
			when "00010110" => data <= '1';
			when "00010111" => data <= '1';
			when "00011000" => data <= '1';
			when "00011001" => data <= '1';
			when "00011010" => data <= '0';
			when "00011011" => data <= '0';
			when "00011100" => data <= '0';
			when "00011101" => data <= '0';
			when "00011110" => data <= '0';
			when "00011111" => data <= '0';
			when "00100000" => data <= '0';
			when "00100001" => data <= '0';
			when "00100010" => data <= '0';
			when "00100011" => data <= '0';
			when "00100100" => data <= '1';
			when "00100101" => data <= '1';
			when "00100110" => data <= '1';
			when "00100111" => data <= '1';
			when "00101000" => data <= '1';
			when "00101001" => data <= '1';
			when "00101010" => data <= '1';
			when "00101011" => data <= '1';
			when "00101100" => data <= '0';
			when "00101101" => data <= '0';
			when "00101110" => data <= '0';
			when "00101111" => data <= '0';
			when "00110000" => data <= '0';
			when "00110001" => data <= '0';
			when "00110010" => data <= '0';
			when "00110011" => data <= '1';
			when "00110100" => data <= '1';
			when "00110101" => data <= '1';
			when "00110110" => data <= '1';
			when "00110111" => data <= '1';
			when "00111000" => data <= '1';
			when "00111001" => data <= '1';
			when "00111010" => data <= '1';
			when "00111011" => data <= '1';
			when "00111100" => data <= '1';
			when "00111101" => data <= '0';
			when "00111110" => data <= '0';
			when "00111111" => data <= '0';
			when "01000000" => data <= '0';
			when "01000001" => data <= '0';
			when "01000010" => data <= '1';
			when "01000011" => data <= '1';
			when "01000100" => data <= '1';
			when "01000101" => data <= '1';
			when "01000110" => data <= '1';
			when "01000111" => data <= '1';
			when "01001000" => data <= '1';
			when "01001001" => data <= '1';
			when "01001010" => data <= '1';
			when "01001011" => data <= '1';
			when "01001100" => data <= '1';
			when "01001101" => data <= '1';
			when "01001110" => data <= '0';
			when "01001111" => data <= '0';
			when "01010000" => data <= '0';
			when "01010001" => data <= '0';
			when "01010010" => data <= '1';
			when "01010011" => data <= '1';
			when "01010100" => data <= '1';
			when "01010101" => data <= '1';
			when "01010110" => data <= '1';
			when "01010111" => data <= '1';
			when "01011000" => data <= '1';
			when "01011001" => data <= '1';
			when "01011010" => data <= '1';
			when "01011011" => data <= '1';
			when "01011100" => data <= '1';
			when "01011101" => data <= '1';
			when "01011110" => data <= '0';
			when "01011111" => data <= '0';
			when "01100000" => data <= '0';
			when "01100001" => data <= '0';
			when "01100010" => data <= '1';
			when "01100011" => data <= '1';
			when "01100100" => data <= '1';
			when "01100101" => data <= '1';
			when "01100110" => data <= '1';
			when "01100111" => data <= '1';
			when "01101000" => data <= '1';
			when "01101001" => data <= '1';
			when "01101010" => data <= '1';
			when "01101011" => data <= '1';
			when "01101100" => data <= '1';
			when "01101101" => data <= '1';
			when "01101110" => data <= '0';
			when "01101111" => data <= '0';
			when "01110000" => data <= '0';
			when "01110001" => data <= '1';
			when "01110010" => data <= '1';
			when "01110011" => data <= '1';
			when "01110100" => data <= '1';
			when "01110101" => data <= '1';
			when "01110110" => data <= '1';
			when "01110111" => data <= '1';
			when "01111000" => data <= '1';
			when "01111001" => data <= '1';
			when "01111010" => data <= '1';
			when "01111011" => data <= '1';
			when "01111100" => data <= '1';
			when "01111101" => data <= '1';
			when "01111110" => data <= '1';
			when "01111111" => data <= '0';
			when "10000000" => data <= '0';
			when "10000001" => data <= '1';
			when "10000010" => data <= '1';
			when "10000011" => data <= '1';
			when "10000100" => data <= '1';
			when "10000101" => data <= '1';
			when "10000110" => data <= '1';
			when "10000111" => data <= '1';
			when "10001000" => data <= '1';
			when "10001001" => data <= '1';
			when "10001010" => data <= '1';
			when "10001011" => data <= '1';
			when "10001100" => data <= '1';
			when "10001101" => data <= '1';
			when "10001110" => data <= '1';
			when "10001111" => data <= '0';
			when "10010000" => data <= '0';
			when "10010001" => data <= '1';
			when "10010010" => data <= '1';
			when "10010011" => data <= '1';
			when "10010100" => data <= '1';
			when "10010101" => data <= '1';
			when "10010110" => data <= '1';
			when "10010111" => data <= '1';
			when "10011000" => data <= '1';
			when "10011001" => data <= '1';
			when "10011010" => data <= '1';
			when "10011011" => data <= '1';
			when "10011100" => data <= '1';
			when "10011101" => data <= '1';
			when "10011110" => data <= '1';
			when "10011111" => data <= '0';
			when "10100000" => data <= '0';
			when "10100001" => data <= '1';
			when "10100010" => data <= '1';
			when "10100011" => data <= '1';
			when "10100100" => data <= '1';
			when "10100101" => data <= '1';
			when "10100110" => data <= '1';
			when "10100111" => data <= '1';
			when "10101000" => data <= '1';
			when "10101001" => data <= '1';
			when "10101010" => data <= '1';
			when "10101011" => data <= '1';
			when "10101100" => data <= '1';
			when "10101101" => data <= '1';
			when "10101110" => data <= '1';
			when "10101111" => data <= '0';
			when "10110000" => data <= '0';
			when "10110001" => data <= '1';
			when "10110010" => data <= '1';
			when "10110011" => data <= '1';
			when "10110100" => data <= '1';
			when "10110101" => data <= '1';
			when "10110110" => data <= '1';
			when "10110111" => data <= '1';
			when "10111000" => data <= '1';
			when "10111001" => data <= '1';
			when "10111010" => data <= '1';
			when "10111011" => data <= '1';
			when "10111100" => data <= '1';
			when "10111101" => data <= '1';
			when "10111110" => data <= '1';
			when "10111111" => data <= '0';
			when "11000000" => data <= '0';
			when "11000001" => data <= '1';
			when "11000010" => data <= '1';
			when "11000011" => data <= '1';
			when "11000100" => data <= '1';
			when "11000101" => data <= '1';
			when "11000110" => data <= '1';
			when "11000111" => data <= '1';
			when "11001000" => data <= '1';
			when "11001001" => data <= '1';
			when "11001010" => data <= '1';
			when "11001011" => data <= '1';
			when "11001100" => data <= '1';
			when "11001101" => data <= '1';
			when "11001110" => data <= '1';
			when "11001111" => data <= '0';
			when "11010000" => data <= '0';
			when "11010001" => data <= '1';
			when "11010010" => data <= '1';
			when "11010011" => data <= '1';
			when "11010100" => data <= '1';
			when "11010101" => data <= '1';
			when "11010110" => data <= '1';
			when "11010111" => data <= '1';
			when "11011000" => data <= '1';
			when "11011001" => data <= '1';
			when "11011010" => data <= '1';
			when "11011011" => data <= '1';
			when "11011100" => data <= '1';
			when "11011101" => data <= '1';
			when "11011110" => data <= '1';
			when "11011111" => data <= '0';
			when "11100000" => data <= '0';
			when "11100001" => data <= '0';
			when "11100010" => data <= '1';
			when "11100011" => data <= '1';
			when "11100100" => data <= '0';
			when "11100101" => data <= '0';
			when "11100110" => data <= '0';
			when "11100111" => data <= '1';
			when "11101000" => data <= '1';
			when "11101001" => data <= '0';
			when "11101010" => data <= '0';
			when "11101011" => data <= '0';
			when "11101100" => data <= '1';
			when "11101101" => data <= '1';
			when "11101110" => data <= '0';
			when "11101111" => data <= '0';
			when "11110000" => data <= '0';
			when "11110001" => data <= '0';
			when "11110010" => data <= '0';
			when "11110011" => data <= '0';
			when "11110100" => data <= '0';
			when "11110101" => data <= '0';
			when "11110110" => data <= '0';
			when "11110111" => data <= '0';
			when "11111000" => data <= '0';
			when "11111001" => data <= '0';
			when "11111010" => data <= '0';
			when "11111011" => data <= '0';
			when "11111100" => data <= '0';
			when "11111101" => data <= '0';
			when "11111110" => data <= '0';
			when "11111111" => data <= '0';
			end case;
		end if;
	end process;
end;