library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity board_map is
  port(
		clk: in std_logic;
		addr : in std_logic_vector(10 downto 0);
		data : out std_logic
  );
end board_map;


architecture synth of board_map is
begin
	process(clk) is begin
		if rising_edge(clk) then
			case addr is
				when "00000000000" => data <= '1';
				when "00000000001" => data <= '1';
				when "00000000010" => data <= '1';
				when "00000000011" => data <= '1';
				when "00000000100" => data <= '1';
				when "00000000101" => data <= '1';
				when "00000000110" => data <= '1';
				when "00000000111" => data <= '1';
				when "00000001000" => data <= '1';
				when "00000001001" => data <= '1';
				when "00000001010" => data <= '1';
				when "00000001011" => data <= '1';
				when "00000001100" => data <= '1';
				when "00000001101" => data <= '1';
				when "00000001110" => data <= '1';
				when "00000001111" => data <= '1';
				when "00000010000" => data <= '1';
				when "00000010001" => data <= '1';
				when "00000010010" => data <= '1';
				when "00000010011" => data <= '1';
				when "00000010100" => data <= '1';
				when "00000010101" => data <= '1';
				when "00000010110" => data <= '1';
				when "00000010111" => data <= '1';
				when "00000011000" => data <= '1';
				when "00000011001" => data <= '1';
				when "00000011010" => data <= '1';
				when "00000011011" => data <= '1';
				when "00000011100" => data <= '1';
				when "00000011101" => data <= '1';
				when "00000011110" => data <= '1';
				when "00000011111" => data <= '1';
				when "00000100000" => data <= '1';
				when "00000100001" => data <= '1';
				when "00000100010" => data <= '1';
				when "00000100011" => data <= '1';
				when "00000100100" => data <= '1';
				when "00000100101" => data <= '1';
				when "00000100110" => data <= '1';
				when "00000100111" => data <= '1';
				when "00000101000" => data <= '1';
				when "00000101001" => data <= '1';
				when "00000101010" => data <= '1';
				when "00000101011" => data <= '1';
				when "00000101100" => data <= '1';
				when "00000101101" => data <= '1';
				when "00000101110" => data <= '1';
				when "00000101111" => data <= '0';
				when "00000110000" => data <= '0';
				when "00000110001" => data <= '0';
				when "00000110010" => data <= '0';
				when "00000110011" => data <= '0';
				when "00000110100" => data <= '0';
				when "00000110101" => data <= '0';
				when "00000110110" => data <= '0';
				when "00000110111" => data <= '0';
				when "00000111000" => data <= '0';
				when "00000111001" => data <= '0';
				when "00000111010" => data <= '0';
				when "00000111011" => data <= '1';
				when "00000111100" => data <= '1';
				when "00000111101" => data <= '0';
				when "00000111110" => data <= '0';
				when "00000111111" => data <= '0';
				when "00001000000" => data <= '0';
				when "00001000001" => data <= '0';
				when "00001000010" => data <= '0';
				when "00001000011" => data <= '0';
				when "00001000100" => data <= '0';
				when "00001000101" => data <= '0';
				when "00001000110" => data <= '0';
				when "00001000111" => data <= '0';
				when "00001001000" => data <= '0';
				when "00001001001" => data <= '1';
				when "00001001010" => data <= '1';
				when "00001001011" => data <= '1';
				when "00001001100" => data <= '1';
				when "00001001101" => data <= '1';
				when "00001001110" => data <= '1';
				when "00001001111" => data <= '1';
				when "00001010000" => data <= '1';
				when "00001010001" => data <= '1';
				when "00001010010" => data <= '1';
				when "00001010011" => data <= '1';
				when "00001010100" => data <= '1';
				when "00001010101" => data <= '1';
				when "00001010110" => data <= '1';
				when "00001010111" => data <= '0';
				when "00001011000" => data <= '1';
				when "00001011001" => data <= '1';
				when "00001011010" => data <= '1';
				when "00001011011" => data <= '1';
				when "00001011100" => data <= '0';
				when "00001011101" => data <= '1';
				when "00001011110" => data <= '1';
				when "00001011111" => data <= '1';
				when "00001100000" => data <= '1';
				when "00001100001" => data <= '1';
				when "00001100010" => data <= '0';
				when "00001100011" => data <= '1';
				when "00001100100" => data <= '1';
				when "00001100101" => data <= '0';
				when "00001100110" => data <= '1';
				when "00001100111" => data <= '1';
				when "00001101000" => data <= '1';
				when "00001101001" => data <= '1';
				when "00001101010" => data <= '1';
				when "00001101011" => data <= '0';
				when "00001101100" => data <= '1';
				when "00001101101" => data <= '1';
				when "00001101110" => data <= '1';
				when "00001101111" => data <= '1';
				when "00001110000" => data <= '0';
				when "00001110001" => data <= '1';
				when "00001110010" => data <= '1';
				when "00001110011" => data <= '1';
				when "00001110100" => data <= '1';
				when "00001110101" => data <= '1';
				when "00001110110" => data <= '1';
				when "00001110111" => data <= '1';
				when "00001111000" => data <= '1';
				when "00001111001" => data <= '1';
				when "00001111010" => data <= '1';
				when "00001111011" => data <= '1';
				when "00001111100" => data <= '1';
				when "00001111101" => data <= '1';
				when "00001111110" => data <= '1';
				when "00001111111" => data <= '0';
				when "00010000000" => data <= '1';
				when "00010000001" => data <= '1';
				when "00010000010" => data <= '1';
				when "00010000011" => data <= '1';
				when "00010000100" => data <= '0';
				when "00010000101" => data <= '1';
				when "00010000110" => data <= '1';
				when "00010000111" => data <= '1';
				when "00010001000" => data <= '1';
				when "00010001001" => data <= '1';
				when "00010001010" => data <= '0';
				when "00010001011" => data <= '1';
				when "00010001100" => data <= '1';
				when "00010001101" => data <= '0';
				when "00010001110" => data <= '1';
				when "00010001111" => data <= '1';
				when "00010010000" => data <= '1';
				when "00010010001" => data <= '1';
				when "00010010010" => data <= '1';
				when "00010010011" => data <= '0';
				when "00010010100" => data <= '1';
				when "00010010101" => data <= '1';
				when "00010010110" => data <= '1';
				when "00010010111" => data <= '1';
				when "00010011000" => data <= '0';
				when "00010011001" => data <= '1';
				when "00010011010" => data <= '1';
				when "00010011011" => data <= '1';
				when "00010011100" => data <= '1';
				when "00010011101" => data <= '1';
				when "00010011110" => data <= '1';
				when "00010011111" => data <= '1';
				when "00010100000" => data <= '1';
				when "00010100001" => data <= '1';
				when "00010100010" => data <= '1';
				when "00010100011" => data <= '1';
				when "00010100100" => data <= '1';
				when "00010100101" => data <= '1';
				when "00010100110" => data <= '1';
				when "00010100111" => data <= '0';
				when "00010101000" => data <= '0';
				when "00010101001" => data <= '0';
				when "00010101010" => data <= '0';
				when "00010101011" => data <= '0';
				when "00010101100" => data <= '0';
				when "00010101101" => data <= '0';
				when "00010101110" => data <= '0';
				when "00010101111" => data <= '0';
				when "00010110000" => data <= '0';
				when "00010110001" => data <= '0';
				when "00010110010" => data <= '0';
				when "00010110011" => data <= '0';
				when "00010110100" => data <= '0';
				when "00010110101" => data <= '0';
				when "00010110110" => data <= '0';
				when "00010110111" => data <= '0';
				when "00010111000" => data <= '0';
				when "00010111001" => data <= '0';
				when "00010111010" => data <= '0';
				when "00010111011" => data <= '0';
				when "00010111100" => data <= '0';
				when "00010111101" => data <= '0';
				when "00010111110" => data <= '0';
				when "00010111111" => data <= '0';
				when "00011000000" => data <= '0';
				when "00011000001" => data <= '1';
				when "00011000010" => data <= '1';
				when "00011000011" => data <= '1';
				when "00011000100" => data <= '1';
				when "00011000101" => data <= '1';
				when "00011000110" => data <= '1';
				when "00011000111" => data <= '1';
				when "00011001000" => data <= '1';
				when "00011001001" => data <= '1';
				when "00011001010" => data <= '1';
				when "00011001011" => data <= '1';
				when "00011001100" => data <= '1';
				when "00011001101" => data <= '1';
				when "00011001110" => data <= '1';
				when "00011001111" => data <= '0';
				when "00011010000" => data <= '1';
				when "00011010001" => data <= '1';
				when "00011010010" => data <= '1';
				when "00011010011" => data <= '1';
				when "00011010100" => data <= '0';
				when "00011010101" => data <= '1';
				when "00011010110" => data <= '1';
				when "00011010111" => data <= '0';
				when "00011011000" => data <= '1';
				when "00011011001" => data <= '1';
				when "00011011010" => data <= '1';
				when "00011011011" => data <= '1';
				when "00011011100" => data <= '1';
				when "00011011101" => data <= '1';
				when "00011011110" => data <= '1';
				when "00011011111" => data <= '1';
				when "00011100000" => data <= '0';
				when "00011100001" => data <= '1';
				when "00011100010" => data <= '1';
				when "00011100011" => data <= '0';
				when "00011100100" => data <= '1';
				when "00011100101" => data <= '1';
				when "00011100110" => data <= '1';
				when "00011100111" => data <= '1';
				when "00011101000" => data <= '0';
				when "00011101001" => data <= '1';
				when "00011101010" => data <= '1';
				when "00011101011" => data <= '1';
				when "00011101100" => data <= '1';
				when "00011101101" => data <= '1';
				when "00011101110" => data <= '1';
				when "00011101111" => data <= '1';
				when "00011110000" => data <= '1';
				when "00011110001" => data <= '1';
				when "00011110010" => data <= '1';
				when "00011110011" => data <= '1';
				when "00011110100" => data <= '1';
				when "00011110101" => data <= '1';
				when "00011110110" => data <= '1';
				when "00011110111" => data <= '0';
				when "00011111000" => data <= '1';
				when "00011111001" => data <= '1';
				when "00011111010" => data <= '1';
				when "00011111011" => data <= '1';
				when "00011111100" => data <= '0';
				when "00011111101" => data <= '1';
				when "00011111110" => data <= '1';
				when "00011111111" => data <= '0';
				when "00100000000" => data <= '1';
				when "00100000001" => data <= '1';
				when "00100000010" => data <= '1';
				when "00100000011" => data <= '1';
				when "00100000100" => data <= '1';
				when "00100000101" => data <= '1';
				when "00100000110" => data <= '1';
				when "00100000111" => data <= '1';
				when "00100001000" => data <= '0';
				when "00100001001" => data <= '1';
				when "00100001010" => data <= '1';
				when "00100001011" => data <= '0';
				when "00100001100" => data <= '1';
				when "00100001101" => data <= '1';
				when "00100001110" => data <= '1';
				when "00100001111" => data <= '1';
				when "00100010000" => data <= '0';
				when "00100010001" => data <= '1';
				when "00100010010" => data <= '1';
				when "00100010011" => data <= '1';
				when "00100010100" => data <= '1';
				when "00100010101" => data <= '1';
				when "00100010110" => data <= '1';
				when "00100010111" => data <= '1';
				when "00100011000" => data <= '1';
				when "00100011001" => data <= '1';
				when "00100011010" => data <= '1';
				when "00100011011" => data <= '1';
				when "00100011100" => data <= '1';
				when "00100011101" => data <= '1';
				when "00100011110" => data <= '1';
				when "00100011111" => data <= '0';
				when "00100100000" => data <= '0';
				when "00100100001" => data <= '0';
				when "00100100010" => data <= '0';
				when "00100100011" => data <= '0';
				when "00100100100" => data <= '0';
				when "00100100101" => data <= '1';
				when "00100100110" => data <= '1';
				when "00100100111" => data <= '0';
				when "00100101000" => data <= '0';
				when "00100101001" => data <= '0';
				when "00100101010" => data <= '0';
				when "00100101011" => data <= '1';
				when "00100101100" => data <= '1';
				when "00100101101" => data <= '0';
				when "00100101110" => data <= '0';
				when "00100101111" => data <= '0';
				when "00100110000" => data <= '0';
				when "00100110001" => data <= '1';
				when "00100110010" => data <= '1';
				when "00100110011" => data <= '0';
				when "00100110100" => data <= '0';
				when "00100110101" => data <= '0';
				when "00100110110" => data <= '0';
				when "00100110111" => data <= '0';
				when "00100111000" => data <= '0';
				when "00100111001" => data <= '1';
				when "00100111010" => data <= '1';
				when "00100111011" => data <= '1';
				when "00100111100" => data <= '1';
				when "00100111101" => data <= '1';
				when "00100111110" => data <= '1';
				when "00100111111" => data <= '1';
				when "00101000000" => data <= '1';
				when "00101000001" => data <= '1';
				when "00101000010" => data <= '1';
				when "00101000011" => data <= '1';
				when "00101000100" => data <= '1';
				when "00101000101" => data <= '1';
				when "00101000110" => data <= '1';
				when "00101000111" => data <= '1';
				when "00101001000" => data <= '1';
				when "00101001001" => data <= '1';
				when "00101001010" => data <= '1';
				when "00101001011" => data <= '1';
				when "00101001100" => data <= '0';
				when "00101001101" => data <= '1';
				when "00101001110" => data <= '1';
				when "00101001111" => data <= '1';
				when "00101010000" => data <= '1';
				when "00101010001" => data <= '1';
				when "00101010010" => data <= '0';
				when "00101010011" => data <= '1';
				when "00101010100" => data <= '1';
				when "00101010101" => data <= '0';
				when "00101010110" => data <= '1';
				when "00101010111" => data <= '1';
				when "00101011000" => data <= '1';
				when "00101011001" => data <= '1';
				when "00101011010" => data <= '1';
				when "00101011011" => data <= '0';
				when "00101011100" => data <= '1';
				when "00101011101" => data <= '1';
				when "00101011110" => data <= '1';
				when "00101011111" => data <= '1';
				when "00101100000" => data <= '1';
				when "00101100001" => data <= '1';
				when "00101100010" => data <= '1';
				when "00101100011" => data <= '1';
				when "00101100100" => data <= '1';
				when "00101100101" => data <= '1';
				when "00101100110" => data <= '1';
				when "00101100111" => data <= '1';
				when "00101101000" => data <= '1';
				when "00101101001" => data <= '1';
				when "00101101010" => data <= '1';
				when "00101101011" => data <= '1';
				when "00101101100" => data <= '1';
				when "00101101101" => data <= '1';
				when "00101101110" => data <= '1';
				when "00101101111" => data <= '1';
				when "00101110000" => data <= '1';
				when "00101110001" => data <= '1';
				when "00101110010" => data <= '1';
				when "00101110011" => data <= '1';
				when "00101110100" => data <= '0';
				when "00101110101" => data <= '1';
				when "00101110110" => data <= '1';
				when "00101110111" => data <= '1';
				when "00101111000" => data <= '1';
				when "00101111001" => data <= '1';
				when "00101111010" => data <= '0';
				when "00101111011" => data <= '1';
				when "00101111100" => data <= '1';
				when "00101111101" => data <= '0';
				when "00101111110" => data <= '1';
				when "00101111111" => data <= '1';
				when "00110000000" => data <= '1';
				when "00110000001" => data <= '1';
				when "00110000010" => data <= '1';
				when "00110000011" => data <= '0';
				when "00110000100" => data <= '1';
				when "00110000101" => data <= '1';
				when "00110000110" => data <= '1';
				when "00110000111" => data <= '1';
				when "00110001000" => data <= '1';
				when "00110001001" => data <= '1';
				when "00110001010" => data <= '1';
				when "00110001011" => data <= '1';
				when "00110001100" => data <= '1';
				when "00110001101" => data <= '1';
				when "00110001110" => data <= '1';
				when "00110001111" => data <= '1';
				when "00110010000" => data <= '1';
				when "00110010001" => data <= '1';
				when "00110010010" => data <= '1';
				when "00110010011" => data <= '1';
				when "00110010100" => data <= '1';
				when "00110010101" => data <= '1';
				when "00110010110" => data <= '1';
				when "00110010111" => data <= '1';
				when "00110011000" => data <= '1';
				when "00110011001" => data <= '1';
				when "00110011010" => data <= '1';
				when "00110011011" => data <= '1';
				when "00110011100" => data <= '0';
				when "00110011101" => data <= '1';
				when "00110011110" => data <= '1';
				when "00110011111" => data <= '0';
				when "00110100000" => data <= '0';
				when "00110100001" => data <= '0';
				when "00110100010" => data <= '0';
				when "00110100011" => data <= '0';
				when "00110100100" => data <= '0';
				when "00110100101" => data <= '0';
				when "00110100110" => data <= '0';
				when "00110100111" => data <= '0';
				when "00110101000" => data <= '0';
				when "00110101001" => data <= '1';
				when "00110101010" => data <= '1';
				when "00110101011" => data <= '0';
				when "00110101100" => data <= '1';
				when "00110101101" => data <= '1';
				when "00110101110" => data <= '1';
				when "00110101111" => data <= '1';
				when "00110110000" => data <= '1';
				when "00110110001" => data <= '1';
				when "00110110010" => data <= '1';
				when "00110110011" => data <= '1';
				when "00110110100" => data <= '1';
				when "00110110101" => data <= '1';
				when "00110110110" => data <= '1';
				when "00110110111" => data <= '1';
				when "00110111000" => data <= '1';
				when "00110111001" => data <= '1';
				when "00110111010" => data <= '1';
				when "00110111011" => data <= '1';
				when "00110111100" => data <= '1';
				when "00110111101" => data <= '1';
				when "00110111110" => data <= '1';
				when "00110111111" => data <= '1';
				when "00111000000" => data <= '1';
				when "00111000001" => data <= '1';
				when "00111000010" => data <= '1';
				when "00111000011" => data <= '1';
				when "00111000100" => data <= '0';
				when "00111000101" => data <= '1';
				when "00111000110" => data <= '1';
				when "00111000111" => data <= '0';
				when "00111001000" => data <= '1';
				when "00111001001" => data <= '1';
				when "00111001010" => data <= '1';
				when "00111001011" => data <= '1';
				when "00111001100" => data <= '1';
				when "00111001101" => data <= '1';
				when "00111001110" => data <= '1';
				when "00111001111" => data <= '1';
				when "00111010000" => data <= '0';
				when "00111010001" => data <= '1';
				when "00111010010" => data <= '1';
				when "00111010011" => data <= '0';
				when "00111010100" => data <= '1';
				when "00111010101" => data <= '1';
				when "00111010110" => data <= '1';
				when "00111010111" => data <= '1';
				when "00111011000" => data <= '1';
				when "00111011001" => data <= '1';
				when "00111011010" => data <= '1';
				when "00111011011" => data <= '1';
				when "00111011100" => data <= '1';
				when "00111011101" => data <= '1';
				when "00111011110" => data <= '1';
				when "00111011111" => data <= '1';
				when "00111100000" => data <= '1';
				when "00111100001" => data <= '1';
				when "00111100010" => data <= '1';
				when "00111100011" => data <= '1';
				when "00111100100" => data <= '1';
				when "00111100101" => data <= '1';
				when "00111100110" => data <= '1';
				when "00111100111" => data <= '1';
				when "00111101000" => data <= '1';
				when "00111101001" => data <= '1';
				when "00111101010" => data <= '1';
				when "00111101011" => data <= '1';
				when "00111101100" => data <= '0';
				when "00111101101" => data <= '1';
				when "00111101110" => data <= '1';
				when "00111101111" => data <= '0';
				when "00111110000" => data <= '1';
				when "00111110001" => data <= '1';
				when "00111110010" => data <= '1';
				when "00111110011" => data <= '1';
				when "00111110100" => data <= '1';
				when "00111110101" => data <= '1';
				when "00111110110" => data <= '1';
				when "00111110111" => data <= '1';
				when "00111111000" => data <= '0';
				when "00111111001" => data <= '1';
				when "00111111010" => data <= '1';
				when "00111111011" => data <= '0';
				when "00111111100" => data <= '1';
				when "00111111101" => data <= '1';
				when "00111111110" => data <= '1';
				when "00111111111" => data <= '1';
				when "01000000000" => data <= '1';
				when "01000000001" => data <= '1';
				when "01000000010" => data <= '1';
				when "01000000011" => data <= '1';
				when "01000000100" => data <= '1';
				when "01000000101" => data <= '1';
				when "01000000110" => data <= '1';
				when "01000000111" => data <= '1';
				when "01000001000" => data <= '1';
				when "01000001001" => data <= '1';
				when "01000001010" => data <= '1';
				when "01000001011" => data <= '1';
				when "01000001100" => data <= '1';
				when "01000001101" => data <= '1';
				when "01000001110" => data <= '0';
				when "01000001111" => data <= '0';
				when "01000010000" => data <= '0';
				when "01000010001" => data <= '0';
				when "01000010010" => data <= '0';
				when "01000010011" => data <= '0';
				when "01000010100" => data <= '0';
				when "01000010101" => data <= '0';
				when "01000010110" => data <= '0';
				when "01000010111" => data <= '0';
				when "01000011000" => data <= '1';
				when "01000011001" => data <= '1';
				when "01000011010" => data <= '1';
				when "01000011011" => data <= '1';
				when "01000011100" => data <= '1';
				when "01000011101" => data <= '1';
				when "01000011110" => data <= '1';
				when "01000011111" => data <= '1';
				when "01000100000" => data <= '0';
				when "01000100001" => data <= '0';
				when "01000100010" => data <= '0';
				when "01000100011" => data <= '0';
				when "01000100100" => data <= '0';
				when "01000100101" => data <= '0';
				when "01000100110" => data <= '0';
				when "01000100111" => data <= '0';
				when "01000101000" => data <= '0';
				when "01000101001" => data <= '0';
				when "01000101010" => data <= '1';
				when "01000101011" => data <= '1';
				when "01000101100" => data <= '1';
				when "01000101101" => data <= '1';
				when "01000101110" => data <= '1';
				when "01000101111" => data <= '1';
				when "01000110000" => data <= '1';
				when "01000110001" => data <= '1';
				when "01000110010" => data <= '1';
				when "01000110011" => data <= '1';
				when "01000110100" => data <= '1';
				when "01000110101" => data <= '1';
				when "01000110110" => data <= '1';
				when "01000110111" => data <= '1';
				when "01000111000" => data <= '1';
				when "01000111001" => data <= '1';
				when "01000111010" => data <= '1';
				when "01000111011" => data <= '1';
				when "01000111100" => data <= '0';
				when "01000111101" => data <= '1';
				when "01000111110" => data <= '1';
				when "01000111111" => data <= '0';
				when "01001000000" => data <= '1';
				when "01001000001" => data <= '1';
				when "01001000010" => data <= '1';
				when "01001000011" => data <= '1';
				when "01001000100" => data <= '1';
				when "01001000101" => data <= '1';
				when "01001000110" => data <= '1';
				when "01001000111" => data <= '1';
				when "01001001000" => data <= '0';
				when "01001001001" => data <= '1';
				when "01001001010" => data <= '1';
				when "01001001011" => data <= '0';
				when "01001001100" => data <= '1';
				when "01001001101" => data <= '1';
				when "01001001110" => data <= '1';
				when "01001001111" => data <= '1';
				when "01001010000" => data <= '1';
				when "01001010001" => data <= '1';
				when "01001010010" => data <= '1';
				when "01001010011" => data <= '1';
				when "01001010100" => data <= '1';
				when "01001010101" => data <= '1';
				when "01001010110" => data <= '1';
				when "01001010111" => data <= '1';
				when "01001011000" => data <= '1';
				when "01001011001" => data <= '1';
				when "01001011010" => data <= '1';
				when "01001011011" => data <= '1';
				when "01001011100" => data <= '1';
				when "01001011101" => data <= '1';
				when "01001011110" => data <= '1';
				when "01001011111" => data <= '1';
				when "01001100000" => data <= '1';
				when "01001100001" => data <= '1';
				when "01001100010" => data <= '1';
				when "01001100011" => data <= '1';
				when "01001100100" => data <= '0';
				when "01001100101" => data <= '1';
				when "01001100110" => data <= '1';
				when "01001100111" => data <= '0';
				when "01001101000" => data <= '1';
				when "01001101001" => data <= '1';
				when "01001101010" => data <= '1';
				when "01001101011" => data <= '1';
				when "01001101100" => data <= '1';
				when "01001101101" => data <= '1';
				when "01001101110" => data <= '1';
				when "01001101111" => data <= '1';
				when "01001110000" => data <= '0';
				when "01001110001" => data <= '1';
				when "01001110010" => data <= '1';
				when "01001110011" => data <= '0';
				when "01001110100" => data <= '1';
				when "01001110101" => data <= '1';
				when "01001110110" => data <= '1';
				when "01001110111" => data <= '1';
				when "01001111000" => data <= '1';
				when "01001111001" => data <= '1';
				when "01001111010" => data <= '1';
				when "01001111011" => data <= '1';
				when "01001111100" => data <= '1';
				when "01001111101" => data <= '1';
				when "01001111110" => data <= '1';
				when "01001111111" => data <= '1';
				when "01010000000" => data <= '1';
				when "01010000001" => data <= '1';
				when "01010000010" => data <= '1';
				when "01010000011" => data <= '1';
				when "01010000100" => data <= '1';
				when "01010000101" => data <= '1';
				when "01010000110" => data <= '1';
				when "01010000111" => data <= '1';
				when "01010001000" => data <= '1';
				when "01010001001" => data <= '1';
				when "01010001010" => data <= '1';
				when "01010001011" => data <= '1';
				when "01010001100" => data <= '0';
				when "01010001101" => data <= '1';
				when "01010001110" => data <= '1';
				when "01010001111" => data <= '0';
				when "01010010000" => data <= '0';
				when "01010010001" => data <= '0';
				when "01010010010" => data <= '0';
				when "01010010011" => data <= '0';
				when "01010010100" => data <= '0';
				when "01010010101" => data <= '0';
				when "01010010110" => data <= '0';
				when "01010010111" => data <= '0';
				when "01010011000" => data <= '0';
				when "01010011001" => data <= '1';
				when "01010011010" => data <= '1';
				when "01010011011" => data <= '0';
				when "01010011100" => data <= '1';
				when "01010011101" => data <= '1';
				when "01010011110" => data <= '1';
				when "01010011111" => data <= '1';
				when "01010100000" => data <= '1';
				when "01010100001" => data <= '1';
				when "01010100010" => data <= '1';
				when "01010100011" => data <= '1';
				when "01010100100" => data <= '1';
				when "01010100101" => data <= '1';
				when "01010100110" => data <= '1';
				when "01010100111" => data <= '1';
				when "01010101000" => data <= '1';
				when "01010101001" => data <= '1';
				when "01010101010" => data <= '1';
				when "01010101011" => data <= '1';
				when "01010101100" => data <= '1';
				when "01010101101" => data <= '1';
				when "01010101110" => data <= '1';
				when "01010101111" => data <= '1';
				when "01010110000" => data <= '1';
				when "01010110001" => data <= '1';
				when "01010110010" => data <= '1';
				when "01010110011" => data <= '1';
				when "01010110100" => data <= '0';
				when "01010110101" => data <= '1';
				when "01010110110" => data <= '1';
				when "01010110111" => data <= '0';
				when "01010111000" => data <= '1';
				when "01010111001" => data <= '1';
				when "01010111010" => data <= '1';
				when "01010111011" => data <= '1';
				when "01010111100" => data <= '1';
				when "01010111101" => data <= '1';
				when "01010111110" => data <= '1';
				when "01010111111" => data <= '1';
				when "01011000000" => data <= '0';
				when "01011000001" => data <= '1';
				when "01011000010" => data <= '1';
				when "01011000011" => data <= '0';
				when "01011000100" => data <= '1';
				when "01011000101" => data <= '1';
				when "01011000110" => data <= '1';
				when "01011000111" => data <= '1';
				when "01011001000" => data <= '1';
				when "01011001001" => data <= '1';
				when "01011001010" => data <= '1';
				when "01011001011" => data <= '1';
				when "01011001100" => data <= '1';
				when "01011001101" => data <= '1';
				when "01011001110" => data <= '1';
				when "01011001111" => data <= '1';
				when "01011010000" => data <= '1';
				when "01011010001" => data <= '1';
				when "01011010010" => data <= '1';
				when "01011010011" => data <= '1';
				when "01011010100" => data <= '1';
				when "01011010101" => data <= '1';
				when "01011010110" => data <= '1';
				when "01011010111" => data <= '1';
				when "01011011000" => data <= '1';
				when "01011011001" => data <= '1';
				when "01011011010" => data <= '1';
				when "01011011011" => data <= '1';
				when "01011011100" => data <= '0';
				when "01011011101" => data <= '1';
				when "01011011110" => data <= '1';
				when "01011011111" => data <= '0';
				when "01011100000" => data <= '1';
				when "01011100001" => data <= '1';
				when "01011100010" => data <= '1';
				when "01011100011" => data <= '1';
				when "01011100100" => data <= '1';
				when "01011100101" => data <= '1';
				when "01011100110" => data <= '1';
				when "01011100111" => data <= '1';
				when "01011101000" => data <= '0';
				when "01011101001" => data <= '1';
				when "01011101010" => data <= '1';
				when "01011101011" => data <= '0';
				when "01011101100" => data <= '1';
				when "01011101101" => data <= '1';
				when "01011101110" => data <= '1';
				when "01011101111" => data <= '1';
				when "01011110000" => data <= '1';
				when "01011110001" => data <= '1';
				when "01011110010" => data <= '1';
				when "01011110011" => data <= '1';
				when "01011110100" => data <= '1';
				when "01011110101" => data <= '1';
				when "01011110110" => data <= '1';
				when "01011110111" => data <= '1';
				when "01011111000" => data <= '1';
				when "01011111001" => data <= '1';
				when "01011111010" => data <= '1';
				when "01011111011" => data <= '1';
				when "01011111100" => data <= '1';
				when "01011111101" => data <= '1';
				when "01011111110" => data <= '1';
				when "01011111111" => data <= '0';
				when "01100000000" => data <= '0';
				when "01100000001" => data <= '0';
				when "01100000010" => data <= '0';
				when "01100000011" => data <= '0';
				when "01100000100" => data <= '0';
				when "01100000101" => data <= '0';
				when "01100000110" => data <= '0';
				when "01100000111" => data <= '0';
				when "01100001000" => data <= '0';
				when "01100001001" => data <= '0';
				when "01100001010" => data <= '0';
				when "01100001011" => data <= '1';
				when "01100001100" => data <= '1';
				when "01100001101" => data <= '0';
				when "01100001110" => data <= '0';
				when "01100001111" => data <= '0';
				when "01100010000" => data <= '0';
				when "01100010001" => data <= '0';
				when "01100010010" => data <= '0';
				when "01100010011" => data <= '0';
				when "01100010100" => data <= '0';
				when "01100010101" => data <= '0';
				when "01100010110" => data <= '0';
				when "01100010111" => data <= '0';
				when "01100011000" => data <= '0';
				when "01100011001" => data <= '1';
				when "01100011010" => data <= '1';
				when "01100011011" => data <= '1';
				when "01100011100" => data <= '1';
				when "01100011101" => data <= '1';
				when "01100011110" => data <= '1';
				when "01100011111" => data <= '1';
				when "01100100000" => data <= '1';
				when "01100100001" => data <= '1';
				when "01100100010" => data <= '1';
				when "01100100011" => data <= '1';
				when "01100100100" => data <= '1';
				when "01100100101" => data <= '1';
				when "01100100110" => data <= '1';
				when "01100100111" => data <= '0';
				when "01100101000" => data <= '1';
				when "01100101001" => data <= '1';
				when "01100101010" => data <= '1';
				when "01100101011" => data <= '1';
				when "01100101100" => data <= '0';
				when "01100101101" => data <= '1';
				when "01100101110" => data <= '1';
				when "01100101111" => data <= '1';
				when "01100110000" => data <= '1';
				when "01100110001" => data <= '1';
				when "01100110010" => data <= '0';
				when "01100110011" => data <= '1';
				when "01100110100" => data <= '1';
				when "01100110101" => data <= '0';
				when "01100110110" => data <= '1';
				when "01100110111" => data <= '1';
				when "01100111000" => data <= '1';
				when "01100111001" => data <= '1';
				when "01100111010" => data <= '1';
				when "01100111011" => data <= '0';
				when "01100111100" => data <= '1';
				when "01100111101" => data <= '1';
				when "01100111110" => data <= '1';
				when "01100111111" => data <= '1';
				when "01101000000" => data <= '0';
				when "01101000001" => data <= '1';
				when "01101000010" => data <= '1';
				when "01101000011" => data <= '1';
				when "01101000100" => data <= '1';
				when "01101000101" => data <= '1';
				when "01101000110" => data <= '1';
				when "01101000111" => data <= '1';
				when "01101001000" => data <= '1';
				when "01101001001" => data <= '1';
				when "01101001010" => data <= '1';
				when "01101001011" => data <= '1';
				when "01101001100" => data <= '1';
				when "01101001101" => data <= '1';
				when "01101001110" => data <= '1';
				when "01101001111" => data <= '0';
				when "01101010000" => data <= '1';
				when "01101010001" => data <= '1';
				when "01101010010" => data <= '1';
				when "01101010011" => data <= '1';
				when "01101010100" => data <= '0';
				when "01101010101" => data <= '1';
				when "01101010110" => data <= '1';
				when "01101010111" => data <= '1';
				when "01101011000" => data <= '1';
				when "01101011001" => data <= '1';
				when "01101011010" => data <= '0';
				when "01101011011" => data <= '1';
				when "01101011100" => data <= '1';
				when "01101011101" => data <= '0';
				when "01101011110" => data <= '1';
				when "01101011111" => data <= '1';
				when "01101100000" => data <= '1';
				when "01101100001" => data <= '1';
				when "01101100010" => data <= '1';
				when "01101100011" => data <= '0';
				when "01101100100" => data <= '1';
				when "01101100101" => data <= '1';
				when "01101100110" => data <= '1';
				when "01101100111" => data <= '1';
				when "01101101000" => data <= '0';
				when "01101101001" => data <= '1';
				when "01101101010" => data <= '1';
				when "01101101011" => data <= '1';
				when "01101101100" => data <= '1';
				when "01101101101" => data <= '1';
				when "01101101110" => data <= '1';
				when "01101101111" => data <= '1';
				when "01101110000" => data <= '1';
				when "01101110001" => data <= '1';
				when "01101110010" => data <= '1';
				when "01101110011" => data <= '1';
				when "01101110100" => data <= '1';
				when "01101110101" => data <= '1';
				when "01101110110" => data <= '1';
				when "01101110111" => data <= '0';
				when "01101111000" => data <= '0';
				when "01101111001" => data <= '0';
				when "01101111010" => data <= '1';
				when "01101111011" => data <= '1';
				when "01101111100" => data <= '0';
				when "01101111101" => data <= '0';
				when "01101111110" => data <= '0';
				when "01101111111" => data <= '0';
				when "01110000000" => data <= '0';
				when "01110000001" => data <= '0';
				when "01110000010" => data <= '0';
				when "01110000011" => data <= '0';
				when "01110000100" => data <= '0';
				when "01110000101" => data <= '0';
				when "01110000110" => data <= '0';
				when "01110000111" => data <= '0';
				when "01110001000" => data <= '0';
				when "01110001001" => data <= '0';
				when "01110001010" => data <= '0';
				when "01110001011" => data <= '0';
				when "01110001100" => data <= '1';
				when "01110001101" => data <= '1';
				when "01110001110" => data <= '0';
				when "01110001111" => data <= '0';
				when "01110010000" => data <= '0';
				when "01110010001" => data <= '1';
				when "01110010010" => data <= '1';
				when "01110010011" => data <= '1';
				when "01110010100" => data <= '1';
				when "01110010101" => data <= '1';
				when "01110010110" => data <= '1';
				when "01110010111" => data <= '1';
				when "01110011000" => data <= '1';
				when "01110011001" => data <= '1';
				when "01110011010" => data <= '1';
				when "01110011011" => data <= '1';
				when "01110011100" => data <= '1';
				when "01110011101" => data <= '1';
				when "01110011110" => data <= '1';
				when "01110011111" => data <= '1';
				when "01110100000" => data <= '1';
				when "01110100001" => data <= '0';
				when "01110100010" => data <= '1';
				when "01110100011" => data <= '1';
				when "01110100100" => data <= '0';
				when "01110100101" => data <= '1';
				when "01110100110" => data <= '1';
				when "01110100111" => data <= '0';
				when "01110101000" => data <= '1';
				when "01110101001" => data <= '1';
				when "01110101010" => data <= '1';
				when "01110101011" => data <= '1';
				when "01110101100" => data <= '1';
				when "01110101101" => data <= '1';
				when "01110101110" => data <= '1';
				when "01110101111" => data <= '1';
				when "01110110000" => data <= '0';
				when "01110110001" => data <= '1';
				when "01110110010" => data <= '1';
				when "01110110011" => data <= '0';
				when "01110110100" => data <= '1';
				when "01110110101" => data <= '1';
				when "01110110110" => data <= '0';
				when "01110110111" => data <= '1';
				when "01110111000" => data <= '1';
				when "01110111001" => data <= '1';
				when "01110111010" => data <= '1';
				when "01110111011" => data <= '1';
				when "01110111100" => data <= '1';
				when "01110111101" => data <= '1';
				when "01110111110" => data <= '1';
				when "01110111111" => data <= '1';
				when "01111000000" => data <= '1';
				when "01111000001" => data <= '1';
				when "01111000010" => data <= '1';
				when "01111000011" => data <= '1';
				when "01111000100" => data <= '1';
				when "01111000101" => data <= '1';
				when "01111000110" => data <= '1';
				when "01111000111" => data <= '1';
				when "01111001000" => data <= '1';
				when "01111001001" => data <= '0';
				when "01111001010" => data <= '1';
				when "01111001011" => data <= '1';
				when "01111001100" => data <= '0';
				when "01111001101" => data <= '1';
				when "01111001110" => data <= '1';
				when "01111001111" => data <= '0';
				when "01111010000" => data <= '1';
				when "01111010001" => data <= '1';
				when "01111010010" => data <= '1';
				when "01111010011" => data <= '1';
				when "01111010100" => data <= '1';
				when "01111010101" => data <= '1';
				when "01111010110" => data <= '1';
				when "01111010111" => data <= '1';
				when "01111011000" => data <= '0';
				when "01111011001" => data <= '1';
				when "01111011010" => data <= '1';
				when "01111011011" => data <= '0';
				when "01111011100" => data <= '1';
				when "01111011101" => data <= '1';
				when "01111011110" => data <= '0';
				when "01111011111" => data <= '1';
				when "01111100000" => data <= '1';
				when "01111100001" => data <= '1';
				when "01111100010" => data <= '1';
				when "01111100011" => data <= '1';
				when "01111100100" => data <= '1';
				when "01111100101" => data <= '1';
				when "01111100110" => data <= '1';
				when "01111100111" => data <= '1';
				when "01111101000" => data <= '1';
				when "01111101001" => data <= '1';
				when "01111101010" => data <= '1';
				when "01111101011" => data <= '1';
				when "01111101100" => data <= '1';
				when "01111101101" => data <= '1';
				when "01111101110" => data <= '1';
				when "01111101111" => data <= '0';
				when "01111110000" => data <= '0';
				when "01111110001" => data <= '0';
				when "01111110010" => data <= '0';
				when "01111110011" => data <= '0';
				when "01111110100" => data <= '0';
				when "01111110101" => data <= '1';
				when "01111110110" => data <= '1';
				when "01111110111" => data <= '0';
				when "01111111000" => data <= '0';
				when "01111111001" => data <= '0';
				when "01111111010" => data <= '0';
				when "01111111011" => data <= '1';
				when "01111111100" => data <= '1';
				when "01111111101" => data <= '0';
				when "01111111110" => data <= '0';
				when "01111111111" => data <= '0';
				when "10000000000" => data <= '0';
				when "10000000001" => data <= '1';
				when "10000000010" => data <= '1';
				when "10000000011" => data <= '0';
				when "10000000100" => data <= '0';
				when "10000000101" => data <= '0';
				when "10000000110" => data <= '0';
				when "10000000111" => data <= '0';
				when "10000001000" => data <= '0';
				when "10000001001" => data <= '1';
				when "10000001010" => data <= '1';
				when "10000001011" => data <= '1';
				when "10000001100" => data <= '1';
				when "10000001101" => data <= '1';
				when "10000001110" => data <= '1';
				when "10000001111" => data <= '1';
				when "10000010000" => data <= '1';
				when "10000010001" => data <= '1';
				when "10000010010" => data <= '1';
				when "10000010011" => data <= '1';
				when "10000010100" => data <= '1';
				when "10000010101" => data <= '1';
				when "10000010110" => data <= '1';
				when "10000010111" => data <= '0';
				when "10000011000" => data <= '1';
				when "10000011001" => data <= '1';
				when "10000011010" => data <= '1';
				when "10000011011" => data <= '1';
				when "10000011100" => data <= '1';
				when "10000011101" => data <= '1';
				when "10000011110" => data <= '1';
				when "10000011111" => data <= '1';
				when "10000100000" => data <= '1';
				when "10000100001" => data <= '1';
				when "10000100010" => data <= '0';
				when "10000100011" => data <= '1';
				when "10000100100" => data <= '1';
				when "10000100101" => data <= '0';
				when "10000100110" => data <= '1';
				when "10000100111" => data <= '1';
				when "10000101000" => data <= '1';
				when "10000101001" => data <= '1';
				when "10000101010" => data <= '1';
				when "10000101011" => data <= '1';
				when "10000101100" => data <= '1';
				when "10000101101" => data <= '1';
				when "10000101110" => data <= '1';
				when "10000101111" => data <= '1';
				when "10000110000" => data <= '0';
				when "10000110001" => data <= '1';
				when "10000110010" => data <= '1';
				when "10000110011" => data <= '1';
				when "10000110100" => data <= '1';
				when "10000110101" => data <= '1';
				when "10000110110" => data <= '1';
				when "10000110111" => data <= '1';
				when "10000111000" => data <= '1';
				when "10000111001" => data <= '1';
				when "10000111010" => data <= '1';
				when "10000111011" => data <= '1';
				when "10000111100" => data <= '1';
				when "10000111101" => data <= '1';
				when "10000111110" => data <= '1';
				when "10000111111" => data <= '0';
				when "10001000000" => data <= '1';
				when "10001000001" => data <= '1';
				when "10001000010" => data <= '1';
				when "10001000011" => data <= '1';
				when "10001000100" => data <= '1';
				when "10001000101" => data <= '1';
				when "10001000110" => data <= '1';
				when "10001000111" => data <= '1';
				when "10001001000" => data <= '1';
				when "10001001001" => data <= '1';
				when "10001001010" => data <= '0';
				when "10001001011" => data <= '1';
				when "10001001100" => data <= '1';
				when "10001001101" => data <= '0';
				when "10001001110" => data <= '1';
				when "10001001111" => data <= '1';
				when "10001010000" => data <= '1';
				when "10001010001" => data <= '1';
				when "10001010010" => data <= '1';
				when "10001010011" => data <= '1';
				when "10001010100" => data <= '1';
				when "10001010101" => data <= '1';
				when "10001010110" => data <= '1';
				when "10001010111" => data <= '1';
				when "10001011000" => data <= '0';
				when "10001011001" => data <= '1';
				when "10001011010" => data <= '1';
				when "10001011011" => data <= '1';
				when "10001011100" => data <= '1';
				when "10001011101" => data <= '1';
				when "10001011110" => data <= '1';
				when "10001011111" => data <= '1';
				when "10001100000" => data <= '1';
				when "10001100001" => data <= '1';
				when "10001100010" => data <= '1';
				when "10001100011" => data <= '1';
				when "10001100100" => data <= '1';
				when "10001100101" => data <= '1';
				when "10001100110" => data <= '1';
				when "10001100111" => data <= '0';
				when "10001101000" => data <= '0';
				when "10001101001" => data <= '0';
				when "10001101010" => data <= '0';
				when "10001101011" => data <= '0';
				when "10001101100" => data <= '0';
				when "10001101101" => data <= '0';
				when "10001101110" => data <= '0';
				when "10001101111" => data <= '0';
				when "10001110000" => data <= '0';
				when "10001110001" => data <= '0';
				when "10001110010" => data <= '0';
				when "10001110011" => data <= '0';
				when "10001110100" => data <= '0';
				when "10001110101" => data <= '0';
				when "10001110110" => data <= '0';
				when "10001110111" => data <= '0';
				when "10001111000" => data <= '0';
				when "10001111001" => data <= '0';
				when "10001111010" => data <= '0';
				when "10001111011" => data <= '0';
				when "10001111100" => data <= '0';
				when "10001111101" => data <= '0';
				when "10001111110" => data <= '0';
				when "10001111111" => data <= '0';
				when "10010000000" => data <= '0';
				when "10010000001" => data <= '1';
				when "10010000010" => data <= '1';
				when "10010000011" => data <= '1';
				when "10010000100" => data <= '1';
				when "10010000101" => data <= '1';
				when "10010000110" => data <= '1';
				when "10010000111" => data <= '1';
				when "10010001000" => data <= '1';
				when "10010001001" => data <= '1';
				when "10010001010" => data <= '1';
				when "10010001011" => data <= '1';
				when "10010001100" => data <= '1';
				when "10010001101" => data <= '1';
				when "10010001110" => data <= '1';
				when "10010001111" => data <= '1';
				when "10010010000" => data <= '1';
				when "10010010001" => data <= '1';
				when "10010010010" => data <= '1';
				when "10010010011" => data <= '1';
				when "10010010100" => data <= '1';
				when "10010010101" => data <= '1';
				when "10010010110" => data <= '1';
				when "10010010111" => data <= '1';
				when "10010011000" => data <= '1';
				when "10010011001" => data <= '1';
				when "10010011010" => data <= '1';
				when "10010011011" => data <= '1';
				when "10010011100" => data <= '1';
				when "10010011101" => data <= '1';
				when "10010011110" => data <= '1';
				when "10010011111" => data <= '1';
				when "10010100000" => data <= '1';
				when "10010100001" => data <= '1';
				when "10010100010" => data <= '1';
				when "10010100011" => data <= '1';
				when "10010100100" => data <= '1';
				when "10010100101" => data <= '1';
				when "10010100110" => data <= '1';
				when "10010100111" => data <= '1';
				when "10010101000" => data <= '1';
				when "10010101001" => data <= '1';
				when "10010101010" => data <= '1';
				when "10010101011" => data <= '1';
				when "10010101100" => data <= '1';
				when "10010101101" => data <= '1';
				when "10010101110" => data <= '1';
				when "10010101111" => data <= '1';
				when others => data <= '0';
			end case;
		end if;
	end process;
end;